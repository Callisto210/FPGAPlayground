library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;
use work.common.all;

entity txcounters is
	port (
		TxClk : in std_logic;
		
		FrameStart : in std_logic;
		FrameSizeOK : out std_logic;
		CurrentField : out txfield_indicator;
		
		IFGStart : in std_logic;
		IFGCntEq12 : out std_logic;
		
		FCSStart : in std_logic;
		FCSCounter : out natural
		
	);
end entity txcounters;

architecture RTL of txcounters is
	--Licznik odpalany jest wraz z rozpoczęciem odbioru adresu MAC
	--Ilość bajtów liczonych musi sie mieścić między 72-1526 bajtów
	--dodatkowo licznik pokazuje część ramki która jest odczytywana
	signal FrameCnt : std_logic_vector(11 downto 0) := (others => '0');
	
	--IFG przy FastEthernet musi odczekać 960 ns czyli 12 bajtów = 96 bitów, 
	--co jest wartością standardową dla ethernet. Dla FE nie przewiduje sie redukcji IFG 
	signal IFGCnt : std_logic_vector(4 downto 0) := (others => '0');
	signal FCSCnt : natural := 0;
	signal IFGCntEq12sig : std_logic;
	
begin	
	IFGCntEq12 <= IFGCntEq12sig;
	FCSCounter <= FCSCnt;
	
	frame_cntr : process (TxClk) is
	begin
		if rising_edge(TxClk) then
			if FrameStart = '0' then
				FrameCnt <= (others => '0');
			elsif FrameStart = '1' then
				FrameCnt <= FrameCnt + 1;
			end if;
		end if;
	end process frame_cntr;
	
	FrameSizeOK <=  '1' when (FrameCnt >= 144 and FrameCnt <= 3052) else
					'0';
								
	CurrentField <= preamble when (FrameCnt >= 0 and FrameCnt < 15) else
					sfd when (FrameCnt >= 15 and FrameCnt < 16) else
					data_pad when (FrameCnt >= 16 and FrameCnt < 136) else
					data;
	
	
	ifg_cntr : process (TxClk) is
	begin
		if rising_edge(TxClk) then
			if IFGStart = '0' then
				IFGCnt <= (others => '0');
			elsif IFGStart = '1' and IFGCntEq12sig = '0' then
				IFGCnt <= IFGCnt + 1;
			end if;
		end if;
	end process ifg_cntr;
	
		IFGCntEq12sig <= '1' when (IFGCnt >= 24) else
					 '0';
	
	fcs_cntr : process (TxClk) is
	begin
		if rising_edge(TxClk) then
			if FCSStart = '0' then
				FCSCnt <= 0;
			elsif FCSStart = '1' then
				FCSCnt <= FCSCnt + 1;
			end if;
		end if;
	end process fcs_cntr;
	
end architecture RTL;
